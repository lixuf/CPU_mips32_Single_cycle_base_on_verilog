module pc_mux1(in0,in1,zero,branch,pc_mux1out);
	input [31:0]in0,in1;
	input zero,branch;
	output [31:0]pc_mux1out;
	assign pc_mux1out=(zero & branch)?in1:in0;
endmodule;